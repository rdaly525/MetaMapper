module mapping_function_3 (
    input data16,
    output O,
    input CLK,
    input ASYNCRESET
);
assign O = data16;
endmodule

