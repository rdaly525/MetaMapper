module coreir_reg_arst #(
    parameter width = 1,
    parameter arst_posedge = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input arst,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg;
  wire real_rst;
  assign real_rst = arst_posedge ? arst : ~arst;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk, posedge real_rst) begin
    if (real_rst) outReg <= init;
    else outReg <= in;
  end
  assign out = outReg;
endmodule

module WrappedPE (
    input [62:0] inst,
    input [15:0] data0,
    input [15:0] data1,
    input bit0,
    input bit1,
    input bit2,
    input clk_en,
    input CLK,
    input ASYNCRESET,
    output [15:0] O0,
    output O1
);
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst18$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst19$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst20$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst21$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst22$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst24$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out;
wire PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_16_eq_inst0_out;
wire [16:0] PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_17_add_inst1_out;
wire [31:0] PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_32_mul_inst0_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out;
wire [7:0] PE_inst0$LUT_inst0$LUT_comb_inst0$magma_Bits_8_and_inst0_out;
wire PE_inst0$PE_comb_inst0$magma_Bit_and_inst0_out;
wire PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out;
wire [1:0] PE_inst0$PE_comb_inst0$self_O0_out_out_out_out;
wire [1:0] PE_inst0$PE_comb_inst0$self_O12_out_out_out_out;
wire [1:0] PE_inst0$PE_comb_inst0$self_O18_out_out_out_out;
wire [1:0] PE_inst0$PE_comb_inst0$self_O24_out_out_out_out;
wire [4:0] PE_inst0$PE_comb_inst0$self_O30_out_out_out_out;
wire [3:0] PE_inst0$PE_comb_inst0$self_O35_out_out_out_out;
wire [1:0] PE_inst0$PE_comb_inst0$self_O6_out_out_out_out;
wire [0:0] PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] PE_inst0$RegisterMode_inst0$Register_inst0$Register_comb_inst0$Mux2xOutUInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] PE_inst0$RegisterMode_inst0$Register_inst0$reg_PR_inst0_out;
wire [0:0] PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] PE_inst0$RegisterMode_inst1$Register_inst0$Register_comb_inst0$Mux2xOutUInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] PE_inst0$RegisterMode_inst1$Register_inst0$reg_PR_inst0_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst2$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out;
wire [0:0] PE_inst0$RegisterMode_inst2$Register_inst0$Register_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst3$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out;
wire [0:0] PE_inst0$RegisterMode_inst3$Register_inst0$Register_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] PE_inst0$RegisterMode_inst4$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out;
wire [0:0] PE_inst0$RegisterMode_inst4$Register_inst0$Register_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out = inst[5] == 1'h1 ? ($signed(PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out)) >= ($signed(PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out)) : PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out >= PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out = inst[5] == 1'h1 ? ($signed(PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out)) <= ($signed(PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out)) : PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out <= PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h03 ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15] : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h05 ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h04 ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0d ? 1'b0 : 1'b0;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0d ? 1'b0 : 1'b0;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0d ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0c ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0c ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst18$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0c ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst19$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0b ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out = inst[5] == 1'h1 ? ($signed(PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out)) >= ($signed(16'h0000)) : PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out >= 16'h0000;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst20$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0b ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst21$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0b ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst18$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst22$coreir_commonlib_mux2x1_inst0$_join_out = (((PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h00) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h01)) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h02)) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h06) ? PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_17_add_inst1_out[16] : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst19$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out = (((PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h00) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h01)) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h02)) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h06) ? ((PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15] & PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15]) & (~ PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_17_add_inst1_out[15])) | (((~ PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15]) & (~ PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15])) & PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_17_add_inst1_out[15]) : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst20$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst24$coreir_commonlib_mux2x1_inst0$_join_out = (((PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h00) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h01)) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h02)) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h06) ? PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_17_add_inst1_out[16] : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst21$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h02) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h06) ? PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0] : 1'b0;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h01 ? 1'b1 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0f ? 1'b0 : 1'b0;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h14 ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h12 ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h13 ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h08 ? 1'b0 : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h01) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h06) ? ~ PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out = (((PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h00) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h01)) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h02)) | (PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h06) ? PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_17_add_inst1_out[15:0] : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0b ? PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_32_mul_inst0_out[15:0] : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0c ? PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_32_mul_inst0_out[23:8] : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0d ? PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_32_mul_inst0_out[31:16] : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h04 ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0] ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h05 ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0] ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h03 ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0] ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out : - PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h08 ? PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0] ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h13 ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out & PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h12 ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out | PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h14 ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out ^ PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$PE_comb_inst0$self_O30_out_out_out_out == 5'h0f ? inst[5] == 1'h1 ? ($signed(PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out)) >>> PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out >> PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out << PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_16_eq_inst0_out = PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out == 16'h0000;
assign PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_17_add_inst1_out = 17'((17'(({1'b0,PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15:0]}) + ({1'b0,PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15:0]}))) + ({1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0]}));
assign PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_32_mul_inst0_out = 32'((inst[5] == 1'h1 ? {PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15:0]} : {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15:0]}) * (inst[5] == 1'h1 ? {PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15],PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15:0]} : {1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,1'b0,PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out[15:0]}));
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out = ((((((((((((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'hf) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h5))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h6))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h7))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h8))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h9))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'ha))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'hb))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'hc))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'hd)) ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst24$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$LUT_inst0$LUT_comb_inst0$magma_Bits_8_and_inst0_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out = (((((((((((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'hd) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h5))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h6))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h7))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h8))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h9))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'ha))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'hb))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'hc)) ? PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_16_eq_inst0_out | (PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out[15] ^ PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out[0]) : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out = ((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3))) ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out[15] : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out = ((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2))) ? ~ PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst22$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out = (((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1)) ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst22$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0)) ? ~ PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_16_eq_inst0_out : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0 ? PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_16_eq_inst0_out : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out = ((((((((((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'hc) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h5))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h6))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h7))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h8))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h9))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'ha))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'hb)) ? (~ PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_16_eq_inst0_out) & (~ (PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out[15] ^ PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out[0])) : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out = (((((((((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'hb) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h5))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h6))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h7))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h8))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h9))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'ha)) ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out[15] ^ PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out = ((((((((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'ha) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h5))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h6))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h7))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h8))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h9)) ? ~ (PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out[15] ^ PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out[0]) : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out = (((((((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h9) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h5))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h6))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h7))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h8)) ? (~ PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst22$coreir_commonlib_mux2x1_inst0$_join_out[0]) | PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_16_eq_inst0_out : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out = ((((((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h8) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h5))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h6))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h7)) ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst22$coreir_commonlib_mux2x1_inst0$_join_out[0] & (~ PE_inst0$ALU_inst0$ALU_comb_inst0$magma_Bits_16_eq_inst0_out) : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out = (((((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h7) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h5))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h6)) ? ~ PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out = ((((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h6) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h5)) ? PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutBit_inst23$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out = (((((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h5) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h0))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h1))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h2)))) & (~ ((PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3) | (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h3)))) & (~ (PE_inst0$PE_comb_inst0$self_O35_out_out_out_out == 4'h4)) ? ~ PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out[15] : PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$LUT_inst0$LUT_comb_inst0$magma_Bits_8_and_inst0_out = (inst[13:6] >> ({1'b0,1'b0,1'b0,1'b0,1'b0,PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0],PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0],PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0]})) & 8'h01;
assign PE_inst0$PE_comb_inst0$magma_Bit_and_inst0_out = (3'h0 == 3'h3) & 1'b0;
assign PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out = (3'h0 == 3'h4) & 1'b0;
assign PE_inst0$PE_comb_inst0$self_O0_out_out_out_out = inst[19:18];
assign PE_inst0$PE_comb_inst0$self_O12_out_out_out_out = inst[55:54];
assign PE_inst0$PE_comb_inst0$self_O18_out_out_out_out = inst[58:57];
assign PE_inst0$PE_comb_inst0$self_O24_out_out_out_out = inst[61:60];
assign PE_inst0$PE_comb_inst0$self_O30_out_out_out_out = inst[4:0];
assign PE_inst0$PE_comb_inst0$self_O35_out_out_out_out = inst[17:14];
assign PE_inst0$PE_comb_inst0$self_O6_out_out_out_out = inst[37:36];
assign PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h3 ? clk_en : 1'b0;
assign PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst0_out ^ 1'b1) ? 1'b1 : PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h0)) ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h0 ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst0_out ^ 1'b1) ? 16'h0000 : PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h3 ? data0 : data0;
assign PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h0 ? inst[35:20] : (PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h0)) ? data0 : ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst0_out ^ 1'b1) ? PE_inst0$RegisterMode_inst0$Register_inst0$reg_PR_inst0_out : PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h3 ? PE_inst0$RegisterMode_inst0$Register_inst0$reg_PR_inst0_out : PE_inst0$RegisterMode_inst0$Register_inst0$reg_PR_inst0_out;
assign PE_inst0$RegisterMode_inst0$Register_inst0$Register_comb_inst0$Mux2xOutUInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out = PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0] ? PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h0 ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out : (PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O0_out_out_out_out == 2'h0)) ? PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$RegisterMode_inst0$RegisterMode_comb_inst0$Mux2xOutUInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$RegisterMode_inst0$Register_inst0$reg_PR_inst0_out;
coreir_reg_arst #(
    .arst_posedge(1'b1),
    .clk_posedge(1'b1),
    .init(16'h0000),
    .width(16)
) PE_inst0$RegisterMode_inst0$Register_inst0$reg_PR_inst0 (
    .clk(CLK),
    .arst(ASYNCRESET),
    .in(PE_inst0$RegisterMode_inst0$Register_inst0$Register_comb_inst0$Mux2xOutUInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .out(PE_inst0$RegisterMode_inst0$Register_inst0$reg_PR_inst0_out)
);
assign PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h3 ? clk_en : 1'b0;
assign PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst0_out ^ 1'b1) ? 1'b1 : PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h0)) ? PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h0 ? PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst0_out ^ 1'b1) ? 16'h0000 : PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h3 ? data1 : data1;
assign PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst8$coreir_commonlib_mux2x16_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h0 ? inst[53:38] : (PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h0)) ? data1 : ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst0_out ^ 1'b1) ? PE_inst0$RegisterMode_inst1$Register_inst0$reg_PR_inst0_out : PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h3 ? PE_inst0$RegisterMode_inst1$Register_inst0$reg_PR_inst0_out : PE_inst0$RegisterMode_inst1$Register_inst0$reg_PR_inst0_out;
assign PE_inst0$RegisterMode_inst1$Register_inst0$Register_comb_inst0$Mux2xOutUInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out = PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0] ? PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h0 ? PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out : (PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O6_out_out_out_out == 2'h0)) ? PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$RegisterMode_inst1$RegisterMode_comb_inst0$Mux2xOutUInt16_inst2$coreir_commonlib_mux2x16_inst0$_join_out : PE_inst0$RegisterMode_inst1$Register_inst0$reg_PR_inst0_out;
coreir_reg_arst #(
    .arst_posedge(1'b1),
    .clk_posedge(1'b1),
    .init(16'h0000),
    .width(16)
) PE_inst0$RegisterMode_inst1$Register_inst0$reg_PR_inst0 (
    .clk(CLK),
    .arst(ASYNCRESET),
    .in(PE_inst0$RegisterMode_inst1$Register_inst0$Register_comb_inst0$Mux2xOutUInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .out(PE_inst0$RegisterMode_inst1$Register_inst0$reg_PR_inst0_out)
);
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h3 ? bit0 : bit0;
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h3 ? clk_en : 1'b0;
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h0 ? PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h0 ? PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h0 ? inst[56] : PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h3 ? PE_inst0$RegisterMode_inst2$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0] : PE_inst0$RegisterMode_inst2$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0];
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out ^ 1'b1) ? 1'b0 : PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out ^ 1'b1) ? 1'b1 : PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out ^ 1'b1) ? PE_inst0$RegisterMode_inst2$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0] : PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h0)) ? PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h0)) ? PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O12_out_out_out_out == 2'h0)) ? bit0 : PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out[0];
coreir_reg_arst #(
    .arst_posedge(1'b1),
    .clk_posedge(1'b1),
    .init(1'h0),
    .width(1)
) PE_inst0$RegisterMode_inst2$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0 (
    .clk(CLK),
    .arst(ASYNCRESET),
    .in(PE_inst0$RegisterMode_inst2$Register_inst0$Register_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .out(PE_inst0$RegisterMode_inst2$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out)
);
assign PE_inst0$RegisterMode_inst2$Register_inst0$Register_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out[0] ? PE_inst0$RegisterMode_inst2$RegisterMode_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst2$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0];
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h3 ? bit1 : bit1;
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h3 ? clk_en : 1'b0;
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h0 ? PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h0 ? PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h0 ? inst[59] : PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h3 ? PE_inst0$RegisterMode_inst3$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0] : PE_inst0$RegisterMode_inst3$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0];
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out ^ 1'b1) ? 1'b0 : PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out ^ 1'b1) ? 1'b1 : PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out ^ 1'b1) ? PE_inst0$RegisterMode_inst3$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0] : PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h0)) ? PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h0)) ? PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O18_out_out_out_out == 2'h0)) ? bit1 : PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out[0];
coreir_reg_arst #(
    .arst_posedge(1'b1),
    .clk_posedge(1'b1),
    .init(1'h0),
    .width(1)
) PE_inst0$RegisterMode_inst3$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0 (
    .clk(CLK),
    .arst(ASYNCRESET),
    .in(PE_inst0$RegisterMode_inst3$Register_inst0$Register_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .out(PE_inst0$RegisterMode_inst3$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out)
);
assign PE_inst0$RegisterMode_inst3$Register_inst0$Register_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out[0] ? PE_inst0$RegisterMode_inst3$RegisterMode_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst3$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0];
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h3 ? bit2 : bit2;
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h3 ? clk_en : 1'b0;
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h0 ? PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h0 ? PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h0 ? inst[62] : PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h3 ? PE_inst0$RegisterMode_inst4$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0] : PE_inst0$RegisterMode_inst4$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0];
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out ^ 1'b1) ? 1'b0 : PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out ^ 1'b1) ? 1'b1 : PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out = ~ (PE_inst0$PE_comb_inst0$magma_Bit_and_inst1_out ^ 1'b1) ? PE_inst0$RegisterMode_inst4$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0] : PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h0)) ? PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h0)) ? PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out = (PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h2) & (~ (PE_inst0$PE_comb_inst0$self_O24_out_out_out_out == 2'h0)) ? bit2 : PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out[0];
coreir_reg_arst #(
    .arst_posedge(1'b1),
    .clk_posedge(1'b1),
    .init(1'h0),
    .width(1)
) PE_inst0$RegisterMode_inst4$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0 (
    .clk(CLK),
    .arst(ASYNCRESET),
    .in(PE_inst0$RegisterMode_inst4$Register_inst0$Register_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .out(PE_inst0$RegisterMode_inst4$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out)
);
assign PE_inst0$RegisterMode_inst4$Register_inst0$Register_comb_inst0$Mux2xOutBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out = PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out[0] ? PE_inst0$RegisterMode_inst4$RegisterMode_comb_inst0$Mux2xOutBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out[0] : PE_inst0$RegisterMode_inst4$Register_inst0$DFF_init0_has_ceFalse_has_resetFalse_has_async_resetTrue_inst0$reg_PR_inst0_out[0];
assign O0 = PE_inst0$ALU_inst0$ALU_comb_inst0$Mux2xOutUInt16_inst17$coreir_commonlib_mux2x16_inst0$_join_out;
assign O1 = PE_inst0$Cond_inst0$Cond_comb_inst0$Mux2xOutBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out[0];
endmodule

